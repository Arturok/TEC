module n_counter #(parameter N= 8)
							(input  logic clk,reset, 
							output logic [N-1:0] q);

always_ff @(posedge clk)
if (reset) q <= 0;
else q <= q + '1;

endmodule